
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;



entity ROM_Array is
    generic(
        N   :   positive :=6; -- number of instructions
        M   :   positive :=32); -- number of bits
    port (
        ADDR:       in STD_LOGIC_VECTOR(N-1 downto 0);
        DATA_OUT:   out STD_LOGIC_VECTOR(M-1 downto 0));
end ROM_Array;


architecture Behavioral of ROM_Array is

    type ROM_array is array (0 to 2**N-1)
        of STD_LOGIC_VECTOR(M-1 downto 0);
         constant ROM    :   ROM_array   := (
        X"e3a0000a", -- asd
        X"e3e01000", -- asd
        X"e3a02002", -- asd
        X"e2802005", -- asd
        X"E2423006", -- asd
        X"E3A0400F", -- asd
        X"E1A050C4", -- asd
        X"E1A06084", -- asd
        X"E5800000", -- asd
        X"E5906000", -- asd
        X"E1550004", -- asd
        X"92809001", -- asd
        X"A280A001", -- asd
        X"e1a00000", -- asd
        X"eb000000", -- asd
        X"e3a0000d", -- asd
        X"eaffffef", -- asd
        X"E2824002", -- asd
        X"e246400d", -- asd
        X"eaffffec", -- asd
        X"00000000",X"00000000",X"00000000",X"00000000",
        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
    );

begin
    DATA_OUT <= ROM(to_integer(unsigned(ADDR)));
end Behavioral;



-- Given Example 
--    constant ROM    :   ROM_array   := (
--        X"E3A00000",X"E3E01000",X"E0812000",X"E24230FF",X"E1A00000",X"EAFFFFF9",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
--    );



--    type ROM_array is array (0 to 2**N-1)
--        of STD_LOGIC_VECTOR(M-1 downto 0);
--            constant ROM    :   ROM_array   := (
--        X"e3a0000a",X"e3e01000",X"e3a02002",X"e2802005",X"e2423006",X"e3a0400f",X"e1a050c4",X"e1a06084",
--        X"E5800000",X"E5906000",X"e1a00000",X"eb000000",X"eafffff2",X"E2824002",X"e246400d",X"eaffffef",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--        X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
--    );
